`include "tx_item.svh"
`include "sequencer.svh"
`include "driver.svh"

module top;
    initial begin
        run_test("run_phase");
    end
endmodule